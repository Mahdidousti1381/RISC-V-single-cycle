module Adder(input [31:0] par_1, input [31:0] par_2, output [31:0] adder_res);
   assign adder_res = par_1 + par_2;
endmodule